module RisingEdge_DFlipFlop(D,clk,Q);
input D; // Data input 
input clk; // clock input 
output Q; // output Q 
always @(posedge clk) 
begin
 Q <= D; 
end 
endmodule 